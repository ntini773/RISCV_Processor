`timescale 1ns/1ps

module NEG_tb;

reg [63:0] A;
wire [63:0] Y;

NEG G1(
    .A(A),
    .Y(Y)
);

initial $monitor("A=%b\nY=%b\n", A, Y);

initial
begin
    $dumpfile("NEG_tb.vcd");
    $dumpvars(0, NEG_tb);

    A = 64'b0000000000000000000000000000000000000000000000000000000000000011; // 3
    #10;

    A = 64'b1111111111111111111111111111111111111111111111111111111111111101; // -3 (in 2's complement)
    #10;

    A = 64'b0000000000000000000000000000000000000000000000000000000000000000; // 0
    #10;

    A = 64'b0000000000000000000000000000000000000000000000000000000000100000; // 32
    #10;

    A = 64'b1111111111111111111111111111111111111111111111111111111111101111; // -33 (in 2's complement)
    #10;

    A = 64'b1111111111111111111111111111111111111111111111111111111111111111; // -1
    #10;

    A = 64'b0000000000000000000000000000000000000000000000000000000000000000; // 0
    #10;

    $finish;
end

endmodule