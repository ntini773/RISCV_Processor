`timescale 1ns/1ps

module OR_tb;

reg [63:0] A;
reg [63:0] B;

wire [63:0] Y;

OR_64 G1(
    .A(A),
    .B(B),
    .Y(Y)
);

initial $monitor("A=%d\nB=%d\nY=%d\n", A, B, Y);

initial
    begin
        $dumpfile("OR_tb.vcd");
        $dumpvars(0, OR_tb);

        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1010101010101010101010101010101010101010101010101010101010101010;
        #10;

        A = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        B = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        #10;

        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;

        A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        B = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        #10;

        A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        B = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        #10;

        A = 64'b1101101101101101101101101101101101101101101101101101101101101101;
        B = 64'b1010101010101010101010101010101010101010101010101010101010101010;
        #10;

        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        #10;

        $finish;
    end

endmodule