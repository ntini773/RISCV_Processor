`timescale 1ns/1ps

module ADD_64_tb;

reg [63:0] A;
reg [63:0] B;
reg Cin;

wire [63:0] S;
wire Cout;
wire Overflow;

ADD_64 UUT(
    .A(A),
    .B(B),
    .Cin(Cin),
    .S(S),
    .Cout(Cout),
    .Overflow(Overflow)
);

initial $monitor("Test case :\nA=%d\nB=%d\nCin=%d\nS=%d\nCout=%d\nOverflow=%d\n", A, B, Cin, S, Cout,Overflow);    

initial
begin
    $dumpfile("ADD_64_tb.vcd");
    $dumpvars(0, ADD_64_tb);

        // Test Case 1: A = 0, B = 0, Cin = 0
        A = 64'b0; B = 64'b0; Cin = 0;
        #10;
        
        // Test Case 2: A = -1, B = -1, Cin = 0
        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        Cin = 0;
        #10;
        
        // Test Case 3: A = 1, B = -1, Cin = 1
        A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        Cin = 1;
        #10;
        
        // Test Case 4: A = 9223372036854775807, B = -1, Cin = 0
        A = 64'b0111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        Cin = 0;
        #10;
        
        // Test Case 5: A = -1, B = -1, Cin = 0
        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        Cin = 0;
        #10;

        // Test Case 6: A = -9223372036854775808, B = -9223372036854775808, Cin = 0
        A = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        B = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        Cin = 0;
        #10;
        
        // Test Case 7: A = 1, B = 1, Cin = 1
        A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        B = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        Cin = 1;
        #10;
        
        // Test Case 8: A = -9223372036854775808, B = -9223372036854775808, Cin = 1
        A = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        B = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        Cin = 1;
        #10

    $finish;
end

endmodule
