`timescale 1ns/1ps

module SUB_64_tb;

reg signed [63:0] A;
reg signed [63:0] B;

wire signed [63:0] S;
wire Overflow;

SUB_64 UUT (
    .a(A),
    .b(B),
    .result(S),
    .Overflow(Overflow)
);

initial $monitor("A=%d\nB=%d\nS=%d\nOverflow=%d\n", A, B, S, Overflow);

initial
begin
        $dumpfile("tb_SUB_64.vcd");
        $dumpvars(0, SUB_64_tb);
        A = 64'b0; B = 64'b0;
        #10;
        
        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;
        
        A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;
        
        A = 64'b0111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;
        
        A = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        #10;

        A = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        B = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        #10;
        
        A = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        B = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        #10;
        
        A = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        B = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        #10

    $finish;
end

endmodule
