`timescale 1ns/1ps

module NOT_64_tb;

reg [63:0] A;

wire [63:0] Y;

NOT_64 UUT (
    .A(A),
    .Y(Y)
);

initial $monitor("A=%b\nY=%b\n", A, Y);

initial
begin
    $dumpfile("NOT_64_tb.vcd");
    $dumpvars(0, NOT_64_tb);

    A = 64'b0000000000000000000000000000000000000000000000000000000000000000; // 0
    #10;

    A = 64'b1111111111111111111111111111111111111111111111111111111111111111; // -1
    #10;

    A = 64'b1000000000000000000000000000000000000000000000000000000000000000; // 2^63
    #10;

    A = 64'b0000000000000000000000001000000000000000000000000000000000000000; // 2^31
    #10;

    A = 64'b0101010101010101010101010101010101010101010101010101010101010101; // Alternating pattern
    #10;

    A = 64'b0000000000000000000000000000000000000000000000000000000000000010; // Only second bit is 1
    #10;

    A = 64'b1100101010011010111001001000110100100000001100111101000011110101; // Random pattern
    #10;

    $finish;
end

endmodule